module fifo
   #(
    parameter DATA_WIDTH=24, // number of bits in a word READ
              ADDR_WIDTH=16  // number of address bits
   )
   (
    input  logic clk, reset,
    input  logic rd, wr,
    input  logic signed [DATA_WIDTH-1:0] w_data,
    output logic empty, full,
    output logic signed [DATA_WIDTH-1:0] r_data
   );

   //signal declaration
   logic [ADDR_WIDTH-1:0] w_addr, r_addr;
   logic wr_en, full_tmp;

   // body
   assign wr_en = wr;
   assign full = full_tmp;
   
   // instantiate fifo control unit
   fifo_ctrl #(.ADDR_WIDTH(ADDR_WIDTH)) c_unit
      (.*, .full(full_tmp));
		
   // instantiate register file
   reg_file 
      #(.DATA_WIDTH(DATA_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) f_unit1 
			(.*);
	

endmodule